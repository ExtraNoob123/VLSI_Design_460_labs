module and_20101021(a, b, c, y);

input a, b, c;
output y; 

and(y, a, b, c);

endmodule 