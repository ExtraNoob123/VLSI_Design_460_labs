module or_20101021(a, b, c, y);

input a, b, c;
output y;

or(y, a, b, c);

endmodule